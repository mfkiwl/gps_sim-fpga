module sat_chan (
    input  logic        clk;
    input  logic[31:0]  freq;
    input  logic[15:0]  gain;
    output logic[15:0]  sout
);

endmodule
